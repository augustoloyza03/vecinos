library verilog;
use verilog.vl_types.all;
entity controlgeneralversion3_4_vlg_vec_tst is
end controlgeneralversion3_4_vlg_vec_tst;
